`timescale 1ns/1ns

module chocorrolTB ();

reg clkTB;

chocorrol choco(.clkIn(clkTB));

always #50 clkTB = ~clkTB;

initial begin
	clkTB = 0;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	#100;
	$stop;
end

endmodule