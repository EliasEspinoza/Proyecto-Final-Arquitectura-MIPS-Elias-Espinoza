`timescale 1ns/1ns

module C_AND (
	input a,
	input b,
	output c
);

assign c = a & b;

endmodule
